`ifndef RKV_WATCHDOG_REG
`define RKV_WATCHDOG_REG

`include "rkv_watchdog_reg.sv"

`endif
