
`ifndef APB_MASTER_SEQUENCER_SV
`define APB_MASTER_SEQUENCER_SV

function apb_master_sequencer::new (string name, uvm_component parent);
  super.new(name, parent);
endfunction : new

`endif // APB_MASTER_SEQUENCER_SV


