`ifndef RKV_WATCHDOG_ELEMENT_SEQUENCES_LIB
`define RKV_WATCHDOG_ELEMENT_SEQUENCES_LIB

`include "rkv_watchdog_base_element_sequence.sv"
`include "rkv_watchdog_inrt_wait_clear.sv"
`include "rkv_watchdog_loadcount.sv"
`include "rkv_watchdog_reg_enable_inrt.sv"
`include "rkv_watchdog_reg_enable_rst.sv"
`include "rkv_watchdog_reg_disable_inrt.sv"
`include "rkv_watchdog_reg_disable_rst.sv"



`endif  // RKV_WATCHDOG_ELEMENT_SEQUENCES_LIB
